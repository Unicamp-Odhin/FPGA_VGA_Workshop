module top (
    input  logic clk, // 50MHz
    input  logic rst_n,

    output logic [7:0] led

);

endmodule
